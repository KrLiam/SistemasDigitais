----------------------------------------------------------------------------------
-- Company:     Federal University of Santa Catarina - UFSC
-- Engineer:    Prof. Dr. Eng. Rafael Luiz Cancian
-- Create Date: 2022
-- Design Name: 
-- Module Name:    registerN
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
-- Dependencies: 
-- Revision: 
-- Revision 1.0 
-- Additional Comments: 
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity RegisterN is
	generic(
		width: positive := 8;
		clearValue: integer := 0
	);
	port(
		-- control
		clock, clear, load: in std_logic;
		-- data
		input: in std_logic_vector(width-1 downto 0);
		output: out std_logic_vector(width-1 downto 0)
	);
end entity;

use ieee.numeric_std.all;

architecture behav0 of RegisterN is
	subtype state is std_logic_vector(width-1 downto 0);
	signal currentState, nextState: state;
begin
	-- next-state logic
	nextState <= std_logic_vector(
			to_unsigned(clearValue, nextState'length)
		) when clear='1' else 
		input when load='1' else 
		currentState;
	
	-- memory element
	
	process(clock) is
	begin
		if rising_edge(clock) then
			currentState <= nextState;
		end if;
	end process;
	
	-- output logic
	output <= currentState;
end architecture;